`timescale 1ns/1ns
module Shifter(dataA, dataB, Signal, dataOut);
    input [31:0] dataA;
    input [4:0] dataB;
    input [2:0] Signal;
    output [31:0] dataOut;

    wire [31:0] one, two, four, eight, sixteen;
    parameter SRL = 3'b011;

    mux2 #(1) box1_1(  1'b0,      dataA[31],  dataB[0], one[31]);
    mux2 #(1) box1_2(  dataA[31], dataA[30],  dataB[0], one[30]);
    mux2 #(1) box1_3(  dataA[30], dataA[29],  dataB[0], one[29]);
    mux2 #(1) box1_4(  dataA[29], dataA[28],  dataB[0], one[28]);
    mux2 #(1) box1_5(  dataA[28], dataA[27],  dataB[0], one[27]);
    mux2 #(1) box1_6(  dataA[27], dataA[26],  dataB[0], one[26]);
    mux2 #(1) box1_7(  dataA[26], dataA[25],  dataB[0], one[25]);
    mux2 #(1) box1_8(  dataA[25], dataA[24],  dataB[0], one[24]);
    mux2 #(1) box1_9(  dataA[24], dataA[23],  dataB[0], one[23]);
    mux2 #(1) box1_10( dataA[23], dataA[22],  dataB[0], one[22]);
    mux2 #(1) box1_11( dataA[22], dataA[21],  dataB[0], one[21]);
    mux2 #(1) box1_12( dataA[21], dataA[20],  dataB[0], one[20]);
    mux2 #(1) box1_13( dataA[20], dataA[19],  dataB[0], one[19]);
    mux2 #(1) box1_14( dataA[19], dataA[18],  dataB[0], one[18]);
    mux2 #(1) box1_15( dataA[18], dataA[17],  dataB[0], one[17]);
    mux2 #(1) box1_16( dataA[17], dataA[16],  dataB[0], one[16]);
    mux2 #(1) box1_17( dataA[16], dataA[15],  dataB[0], one[15]);
    mux2 #(1) box1_18( dataA[15], dataA[14],  dataB[0], one[14]);
    mux2 #(1) box1_19( dataA[14], dataA[13],  dataB[0], one[13]);
    mux2 #(1) box1_20( dataA[13], dataA[12],  dataB[0], one[12]);
    mux2 #(1) box1_21( dataA[12], dataA[11],  dataB[0], one[11]);
    mux2 #(1) box1_22( dataA[11], dataA[10],  dataB[0], one[10]);
    mux2 #(1) box1_23( dataA[10], dataA[9],   dataB[0], one[9]);
    mux2 #(1) box1_24( dataA[9],  dataA[8],   dataB[0], one[8]);
    mux2 #(1) box1_25( dataA[8],  dataA[7],   dataB[0], one[7]);
    mux2 #(1) box1_26( dataA[7],  dataA[6],   dataB[0], one[6]);
    mux2 #(1) box1_27( dataA[6],  dataA[5],   dataB[0], one[5]);
    mux2 #(1) box1_28( dataA[5],  dataA[4],   dataB[0], one[4]);
    mux2 #(1) box1_29( dataA[4],  dataA[3],   dataB[0], one[3]);
    mux2 #(1) box1_30( dataA[3],  dataA[2],   dataB[0], one[2]);
    mux2 #(1) box1_31( dataA[2],  dataA[1],   dataB[0], one[1]);
    mux2 #(1) box1_32( dataA[1],  dataA[0],   dataB[0], one[0]);


    mux2 #(1) box2_1(  1'b0,    one[31],  dataB[1], two[31]);
    mux2 #(1) box2_2(  1'b0,    one[30],  dataB[1], two[30]);
    mux2 #(1) box2_3(  one[31], one[29],  dataB[1], two[29]);
    mux2 #(1) box2_4(  one[30], one[28],  dataB[1], two[28]);
    mux2 #(1) box2_5(  one[29], one[27],  dataB[1], two[27]);
    mux2 #(1) box2_6(  one[28], one[26],  dataB[1], two[26]);
    mux2 #(1) box2_7(  one[27], one[25],  dataB[1], two[25]);
    mux2 #(1) box2_8(  one[26], one[24],  dataB[1], two[24]);
    mux2 #(1) box2_9(  one[25], one[23],  dataB[1], two[23]);
    mux2 #(1) box2_10( one[24], one[22],  dataB[1], two[22]);
    mux2 #(1) box2_11( one[23], one[21],  dataB[1], two[21]);
    mux2 #(1) box2_12( one[22], one[20],  dataB[1], two[20]);
    mux2 #(1) box2_13( one[21], one[19],  dataB[1], two[19]);
    mux2 #(1) box2_14( one[20], one[18],  dataB[1], two[18]); 
    mux2 #(1) box2_15( one[19], one[17],  dataB[1], two[17]);
    mux2 #(1) box2_16( one[18], one[16],  dataB[1], two[16]);
    mux2 #(1) box2_17( one[17], one[15],  dataB[1], two[15]);
    mux2 #(1) box2_18( one[16], one[14],  dataB[1], two[14]);
    mux2 #(1) box2_19( one[15], one[13],  dataB[1], two[13]);
    mux2 #(1) box2_20( one[14], one[12],  dataB[1], two[12]);
    mux2 #(1) box2_21( one[13], one[11],  dataB[1], two[11]);
    mux2 #(1) box2_22( one[12], one[10],  dataB[1], two[10]);
    mux2 #(1) box2_23( one[11], one[9],   dataB[1], two[9]);
    mux2 #(1) box2_24( one[10], one[8],   dataB[1], two[8]);
    mux2 #(1) box2_25( one[9],  one[7],   dataB[1], two[7]);
    mux2 #(1) box2_26( one[8],  one[6],   dataB[1], two[6]);
    mux2 #(1) box2_27( one[7],  one[5],   dataB[1], two[5]);
    mux2 #(1) box2_28( one[6],  one[4],   dataB[1], two[4]);
    mux2 #(1) box2_29( one[5],  one[3],   dataB[1], two[3]);
    mux2 #(1) box2_30( one[4],  one[2],   dataB[1], two[2]);
    mux2 #(1) box2_31( one[3],  one[1],   dataB[1], two[1]);
    mux2 #(1) box2_32( one[2],  one[0],   dataB[1], two[0]);


    mux2 #(1) box3_1(  1'b0,    two[31],  dataB[2], four[31]);
    mux2 #(1) box3_2(  1'b0,    two[30],  dataB[2], four[30]);
    mux2 #(1) box3_3(  1'b0,    two[29],  dataB[2], four[29]);
    mux2 #(1) box3_4(  1'b0,    two[28],  dataB[2], four[28]);
    mux2 #(1) box3_5(  two[31], two[27],  dataB[2], four[27]);
    mux2 #(1) box3_6(  two[30], two[26],  dataB[2], four[26]);
    mux2 #(1) box3_7(  two[29], two[25],  dataB[2], four[25]);
    mux2 #(1) box3_8(  two[28], two[24],  dataB[2], four[24]);
    mux2 #(1) box3_9(  two[27], two[23],  dataB[2], four[23]);
    mux2 #(1) box3_10( two[26], two[22],  dataB[2], four[22]);
    mux2 #(1) box3_11( two[25], two[21],  dataB[2], four[21]);
    mux2 #(1) box3_12( two[24], two[20],  dataB[2], four[20]);
    mux2 #(1) box3_13( two[23], two[19],  dataB[2], four[19]);
    mux2 #(1) box3_14( two[22], two[18],  dataB[2], four[18]);
    mux2 #(1) box3_15( two[21], two[17],  dataB[2], four[17]);
    mux2 #(1) box3_16( two[20], two[16],  dataB[2], four[16]);
    mux2 #(1) box3_17( two[19], two[15],  dataB[2], four[15]);
    mux2 #(1) box3_18( two[18], two[14],  dataB[2], four[14]);
    mux2 #(1) box3_19( two[17], two[13],  dataB[2], four[13]);
    mux2 #(1) box3_20( two[16], two[12],  dataB[2], four[12]);
    mux2 #(1) box3_21( two[15], two[11],  dataB[2], four[11]);
    mux2 #(1) box3_22( two[14], two[10],  dataB[2], four[10]);
    mux2 #(1) box3_23( two[13], two[9],   dataB[2], four[9]);
    mux2 #(1) box3_24( two[12], two[8],   dataB[2], four[8]);
    mux2 #(1) box3_25( two[11], two[7],   dataB[2], four[7]);
    mux2 #(1) box3_26( two[10], two[6],   dataB[2], four[6]);
    mux2 #(1) box3_27( two[9],  two[5],   dataB[2], four[5]);
    mux2 #(1) box3_28( two[8],  two[4],   dataB[2], four[4]);
    mux2 #(1) box3_29( two[7],  two[3],   dataB[2], four[3]);
    mux2 #(1) box3_30( two[6],  two[2],   dataB[2], four[2]);
    mux2 #(1) box3_31( two[5],  two[1],   dataB[2], four[1]);
    mux2 #(1) box3_32( two[4],  two[0],   dataB[2], four[0]);


    mux2 #(1) box4_1(  1'b0,     four[31],  dataB[3], eight[31]);
    mux2 #(1) box4_2(  1'b0,     four[30],  dataB[3], eight[30]);
    mux2 #(1) box4_3(  1'b0,     four[29],  dataB[3], eight[29]);
    mux2 #(1) box4_4(  1'b0,     four[28],  dataB[3], eight[28]);
    mux2 #(1) box4_5(  1'b0,     four[27],  dataB[3], eight[27]);
    mux2 #(1) box4_6(  1'b0,     four[26],  dataB[3], eight[26]);
    mux2 #(1) box4_7(  1'b0,     four[25],  dataB[3], eight[25]);
    mux2 #(1) box4_8(  1'b0,     four[24],  dataB[3], eight[24]);
    mux2 #(1) box4_9(  four[31], four[23],  dataB[3], eight[23]);
    mux2 #(1) box4_10( four[30], four[22],  dataB[3], eight[22]);
    mux2 #(1) box4_11( four[29], four[21],  dataB[3], eight[21]);
    mux2 #(1) box4_12( four[28], four[20],  dataB[3], eight[20]);
    mux2 #(1) box4_13( four[27], four[19],  dataB[3], eight[19]);
    mux2 #(1) box4_14( four[26], four[18],  dataB[3], eight[18]);
    mux2 #(1) box4_15( four[25], four[17],  dataB[3], eight[17]);
    mux2 #(1) box4_16( four[24], four[16],  dataB[3], eight[16]);
    mux2 #(1) box4_17( four[23], four[15],  dataB[3], eight[15]);
    mux2 #(1) box4_18( four[22], four[14],  dataB[3], eight[14]);
    mux2 #(1) box4_19( four[21], four[13],  dataB[3], eight[13]);
    mux2 #(1) box4_20( four[20], four[12],  dataB[3], eight[12]);
    mux2 #(1) box4_21( four[19], four[11],  dataB[3], eight[11]);
    mux2 #(1) box4_22( four[18], four[10],  dataB[3], eight[10]);
    mux2 #(1) box4_23( four[17], four[9],   dataB[3], eight[9]);
    mux2 #(1) box4_24( four[16], four[8],   dataB[3], eight[8]);
    mux2 #(1) box4_25( four[15], four[7],   dataB[3], eight[7]);
    mux2 #(1) box4_26( four[14], four[6],   dataB[3], eight[6]);
    mux2 #(1) box4_27( four[13], four[5],   dataB[3], eight[5]);
    mux2 #(1) box4_28( four[12], four[4],   dataB[3], eight[4]);
    mux2 #(1) box4_29( four[11], four[3],   dataB[3], eight[3]);
    mux2 #(1) box4_30( four[10], four[2],   dataB[3], eight[2]);
    mux2 #(1) box4_31( four[9],  four[1],   dataB[3], eight[1]);
    mux2 #(1) box4_32( four[8],  four[0],   dataB[3], eight[0]);


    mux2 #(1) box5_1(  1'b0,      eight[31], dataB[4], sixteen[31]);
    mux2 #(1) box5_2(  1'b0,      eight[30], dataB[4], sixteen[30]);
    mux2 #(1) box5_3(  1'b0,      eight[29], dataB[4], sixteen[29]);
    mux2 #(1) box5_4(  1'b0,      eight[28], dataB[4], sixteen[28]);
    mux2 #(1) box5_5(  1'b0,      eight[27], dataB[4], sixteen[27]);
    mux2 #(1) box5_6(  1'b0,      eight[26], dataB[4], sixteen[26]);
    mux2 #(1) box5_7(  1'b0,      eight[25], dataB[4], sixteen[25]);
    mux2 #(1) box5_8(  1'b0,      eight[24], dataB[4], sixteen[24]);
    mux2 #(1) box5_9(  1'b0,      eight[23], dataB[4], sixteen[23]);
    mux2 #(1) box5_10( 1'b0,      eight[22], dataB[4], sixteen[22]);
    mux2 #(1) box5_11( 1'b0,      eight[21], dataB[4], sixteen[21]);
    mux2 #(1) box5_12( 1'b0,      eight[20], dataB[4], sixteen[20]);
    mux2 #(1) box5_13( 1'b0,      eight[19], dataB[4], sixteen[19]);
    mux2 #(1) box5_14( 1'b0,      eight[18], dataB[4], sixteen[18]);
    mux2 #(1) box5_15( 1'b0,      eight[17], dataB[4], sixteen[17]);
    mux2 #(1) box5_16( 1'b0,      eight[16], dataB[4], sixteen[16]);
    mux2 #(1) box5_17( eight[31], eight[15], dataB[4], sixteen[15]);
    mux2 #(1) box5_18( eight[30], eight[14], dataB[4], sixteen[14]);
    mux2 #(1) box5_19( eight[29], eight[13], dataB[4], sixteen[13]);
    mux2 #(1) box5_20( eight[28], eight[12], dataB[4], sixteen[12]);
    mux2 #(1) box5_21( eight[27], eight[11], dataB[4], sixteen[11]);
    mux2 #(1) box5_22( eight[26], eight[10], dataB[4], sixteen[10]);
    mux2 #(1) box5_23( eight[25], eight[9],  dataB[4], sixteen[9]);
    mux2 #(1) box5_24( eight[24], eight[8],  dataB[4], sixteen[8]);
    mux2 #(1) box5_25( eight[23], eight[7],  dataB[4], sixteen[7]);
    mux2 #(1) box5_26( eight[22], eight[6],  dataB[4], sixteen[6]);
    mux2 #(1) box5_27( eight[21], eight[5],  dataB[4], sixteen[5]);
    mux2 #(1) box5_28( eight[20], eight[4],  dataB[4], sixteen[4]);
    mux2 #(1) box5_29( eight[19], eight[3],  dataB[4], sixteen[3]);
    mux2 #(1) box5_30( eight[18], eight[2],  dataB[4], sixteen[2]);
    mux2 #(1) box5_31( eight[17], eight[1],  dataB[4], sixteen[1]);
    mux2 #(1) box5_32( eight[16], eight[0],  dataB[4], sixteen[0]);
    
    assign dataOut = Signal == SRL ? sixteen : 32'b0;
endmodule